`timescale 1ns / 1ps

module top_hardware_accelerator #(parameter Width = 32) 
(	input clk,
	input reset_n,
	input write,
	input read,
	input [8:0] address,
	input [31:0] writedata,
	output wire OutInt,
	output wire[31:0] readdata);

	wire [Width-1:0] A11InReal,A11InImag,A12InReal,A12InImag,A13InReal,A13InImag,A14InReal,A14InImag,
		B11InReal,B11InImag,B21InReal,B21InImag,B31InReal,B31InImag,B41InReal,B41InImag,
		A21InReal,A21InImag,A22InReal,A22InImag,A23InReal,A23InImag,A24InReal,A24InImag,
		B12InReal,B12InImag,B22InReal,B22InImag,B32InReal,B32InImag,B42InReal,B42InImag,
		A31InReal,A31InImag,A32InReal,A32InImag,A33InReal,A33InImag,A34InReal,A34InImag,
		B13InReal,B13InImag,B23InReal,B23InImag,B33InReal,B33InImag,B43InReal,B43InImag,
		A41InReal,A41InImag,A42InReal,A42InImag,A43InReal,A43InImag,A44InReal,A44InImag,
		B14InReal,B14InImag,B24InReal,B24InImag,B34InReal,B34InImag,B44InReal,B44InImag;
		
	wire [Width-1:0] Out11Real,Out11Imag,Out12Real,Out12Imag,Out13Real,Out13Imag,Out14Real,Out14Imag,
		Out21Real,Out21Imag,Out22Real,Out22Imag,Out23Real,Out23Imag,Out24Real,Out24Imag,
		Out31Real,Out31Imag,Out32Real,Out32Imag,Out33Real,Out33Imag,Out34Real,Out34Imag,
		Out41Real,Out41Imag,Out42Real,Out42Imag,Out43Real,Out43Imag,Out44Real,Out44Imag;
		
	wire EnableListo,Error,Start;
	
	MultiplicadorMatrices #(.Width(Width)) MultiplicadorMatricescopia (
    .CLK(clk), 
    .Enable(1'b1), 
    .MasterReset(~reset_n), ///////////////////////////
    .Start(Start), 
    .A11InReal(A11InReal), 
    .A11InImag(A11InImag), 
    .A12InReal(A12InReal), 
    .A12InImag(A12InImag), 
    .A13InReal(A13InReal), 
    .A13InImag(A13InImag), 
    .A14InReal(A14InReal), 
    .A14InImag(A14InImag), 
    .B11InReal(B11InReal), 
    .B11InImag(B11InImag), 
    .B21InReal(B21InReal), 
    .B21InImag(B21InImag), 
    .B31InReal(B31InReal), 
    .B31InImag(B31InImag), 
    .B41InReal(B41InReal), 
    .B41InImag(B41InImag), 
    .A21InReal(A21InReal), 
    .A21InImag(A21InImag), 
    .A22InReal(A22InReal), 
    .A22InImag(A22InImag), 
    .A23InReal(A23InReal), 
    .A23InImag(A23InImag), 
    .A24InReal(A24InReal), 
    .A24InImag(A24InImag), 
    .B12InReal(B12InReal), 
    .B12InImag(B12InImag), 
    .B22InReal(B22InReal), 
    .B22InImag(B22InImag), 
    .B32InReal(B32InReal), 
    .B32InImag(B32InImag), 
    .B42InReal(B42InReal), 
    .B42InImag(B42InImag), 
    .A31InReal(A31InReal), 
    .A31InImag(A31InImag), 
    .A32InReal(A32InReal), 
    .A32InImag(A32InImag), 
    .A33InReal(A33InReal), 
    .A33InImag(A33InImag), 
    .A34InReal(A34InReal), 
    .A34InImag(A34InImag), 
    .B13InReal(B13InReal), 
    .B13InImag(B13InImag), 
    .B23InReal(B23InReal), 
    .B23InImag(B23InImag), 
    .B33InReal(B33InReal), 
    .B33InImag(B33InImag), 
    .B43InReal(B43InReal), 
    .B43InImag(B43InImag), 
    .A41InReal(A41InReal), 
    .A41InImag(A41InImag), 
    .A42InReal(A42InReal), 
    .A42InImag(A42InImag), 
    .A43InReal(A43InReal), 
    .A43InImag(A43InImag), 
    .A44InReal(A44InReal), 
    .A44InImag(A44InImag), 
    .B14InReal(B14InReal), 
    .B14InImag(B14InImag), 
    .B24InReal(B24InReal), 
    .B24InImag(B24InImag), 
    .B34InReal(B34InReal), 
    .B34InImag(B34InImag), 
    .B44InReal(B44InReal), 
    .B44InImag(B44InImag), 
    .Out11Real(Out11Real), 
    .Out11Imag(Out11Imag), 
    .Out12Real(Out12Real), 
    .Out12Imag(Out12Imag), 
    .Out13Real(Out13Real), 
    .Out13Imag(Out13Imag), 
    .Out14Real(Out14Real), 
    .Out14Imag(Out14Imag), 
    .Out21Real(Out21Real), 
    .Out21Imag(Out21Imag), 
    .Out22Real(Out22Real), 
    .Out22Imag(Out22Imag), 
    .Out23Real(Out23Real), 
    .Out23Imag(Out23Imag), 
    .Out24Real(Out24Real), 
    .Out24Imag(Out24Imag), 
    .Out31Real(Out31Real), 
    .Out31Imag(Out31Imag), 
    .Out32Real(Out32Real), 
    .Out32Imag(Out32Imag), 
    .Out33Real(Out33Real), 
    .Out33Imag(Out33Imag), 
    .Out34Real(Out34Real), 
    .Out34Imag(Out34Imag), 
    .Out41Real(Out41Real), 
    .Out41Imag(Out41Imag), 
    .Out42Real(Out42Real), 
    .Out42Imag(Out42Imag), 
    .Out43Real(Out43Real), 
    .Out43Imag(Out43Imag), 
    .Out44Real(Out44Real), 
    .Out44Imag(Out44Imag), 
    .Listo(EnableListo), 
    .Error(Error)
    );

	// Instantiate the module
	RegistroLoad #(.Width(Width)) RegistroLoadcopia (
    .CLK(clk), 
    .MasterReset(~reset_n | EnableListo), 
    .InDatos(writedata), 
    .Write(write), 
    .Address(address), 
    .A11InReal(A11InReal), 
    .A11InImag(A11InImag), 
    .A12InReal(A12InReal), 
    .A12InImag(A12InImag), 
    .A13InReal(A13InReal), 
    .A13InImag(A13InImag), 
    .A14InReal(A14InReal), 
    .A14InImag(A14InImag), 
    .B11InReal(B11InReal), 
    .B11InImag(B11InImag), 
    .B21InReal(B21InReal), 
    .B21InImag(B21InImag), 
    .B31InReal(B31InReal), 
    .B31InImag(B31InImag), 
    .B41InReal(B41InReal), 
    .B41InImag(B41InImag), 
    .A21InReal(A21InReal), 
    .A21InImag(A21InImag), 
    .A22InReal(A22InReal), 
    .A22InImag(A22InImag), 
    .A23InReal(A23InReal), 
    .A23InImag(A23InImag), 
    .A24InReal(A24InReal), 
    .A24InImag(A24InImag), 
    .B12InReal(B12InReal), 
    .B12InImag(B12InImag), 
    .B22InReal(B22InReal), 
    .B22InImag(B22InImag), 
    .B32InReal(B32InReal), 
    .B32InImag(B32InImag), 
    .B42InReal(B42InReal), 
    .B42InImag(B42InImag), 
    .A31InReal(A31InReal), 
    .A31InImag(A31InImag), 
    .A32InReal(A32InReal), 
    .A32InImag(A32InImag), 
    .A33InReal(A33InReal), 
    .A33InImag(A33InImag), 
    .A34InReal(A34InReal), 
    .A34InImag(A34InImag), 
    .B13InReal(B13InReal), 
    .B13InImag(B13InImag), 
    .B23InReal(B23InReal), 
    .B23InImag(B23InImag), 
    .B33InReal(B33InReal), 
    .B33InImag(B33InImag), 
    .B43InReal(B43InReal), 
    .B43InImag(B43InImag), 
    .A41InReal(A41InReal), 
    .A41InImag(A41InImag), 
    .A42InReal(A42InReal), 
    .A42InImag(A42InImag), 
    .A43InReal(A43InReal), 
    .A43InImag(A43InImag), 
    .A44InReal(A44InReal), 
    .A44InImag(A44InImag), 
    .B14InReal(B14InReal), 
    .B14InImag(B14InImag), 
    .B24InReal(B24InReal), 
    .B24InImag(B24InImag), 
    .B34InReal(B34InReal), 
    .B34InImag(B34InImag), 
    .B44InReal(B44InReal), 
    .B44InImag(B44InImag), 
    .Start(Start)
    );

	
	// Instantiate the module
	MuxSalida #(.Width(Width)) MuxSalidacopia (
    .Read(read), 
    .Address(address), 
	 .A11InReal(A11InReal), 
    .A11InImag(A11InImag), 
    .A12InReal(A12InReal), 
    .A12InImag(A12InImag), 
    .A13InReal(A13InReal), 
    .A13InImag(A13InImag), 
    .A14InReal(A14InReal), 
    .A14InImag(A14InImag), 
    .B11InReal(B11InReal), 
    .B11InImag(B11InImag), 
    .B21InReal(B21InReal), 
    .B21InImag(B21InImag), 
    .B31InReal(B31InReal), 
    .B31InImag(B31InImag), 
    .B41InReal(B41InReal), 
    .B41InImag(B41InImag), 
    .A21InReal(A21InReal), 
    .A21InImag(A21InImag), 
    .A22InReal(A22InReal), 
    .A22InImag(A22InImag), 
    .A23InReal(A23InReal), 
    .A23InImag(A23InImag), 
    .A24InReal(A24InReal), 
    .A24InImag(A24InImag), 
    .B12InReal(B12InReal), 
    .B12InImag(B12InImag), 
    .B22InReal(B22InReal), 
    .B22InImag(B22InImag), 
    .B32InReal(B32InReal), 
    .B32InImag(B32InImag), 
    .B42InReal(B42InReal), 
    .B42InImag(B42InImag), 
    .A31InReal(A31InReal), 
    .A31InImag(A31InImag), 
    .A32InReal(A32InReal), 
    .A32InImag(A32InImag), 
    .A33InReal(A33InReal), 
    .A33InImag(A33InImag), 
    .A34InReal(A34InReal), 
    .A34InImag(A34InImag), 
    .B13InReal(B13InReal), 
    .B13InImag(B13InImag), 
    .B23InReal(B23InReal), 
    .B23InImag(B23InImag), 
    .B33InReal(B33InReal), 
    .B33InImag(B33InImag), 
    .B43InReal(B43InReal), 
    .B43InImag(B43InImag), 
    .A41InReal(A41InReal), 
    .A41InImag(A41InImag), 
    .A42InReal(A42InReal), 
    .A42InImag(A42InImag), 
    .A43InReal(A43InReal), 
    .A43InImag(A43InImag), 
    .A44InReal(A44InReal), 
    .A44InImag(A44InImag), 
    .B14InReal(B14InReal), 
    .B14InImag(B14InImag), 
    .B24InReal(B24InReal), 
    .B24InImag(B24InImag), 
    .B34InReal(B34InReal), 
    .B34InImag(B34InImag), 
    .B44InReal(B44InReal), 
    .B44InImag(B44InImag), 
	 .Start(Start),
	 
    .Out11Real(Out11Real), 
    .Out11Imag(Out11Imag), 
    .Out12Real(Out12Real), 
    .Out12Imag(Out12Imag), 
    .Out13Real(Out13Real), 
    .Out13Imag(Out13Imag), 
    .Out14Real(Out14Real), 
    .Out14Imag(Out14Imag), 
    .Out21Real(Out21Real), 
    .Out21Imag(Out21Imag), 
    .Out22Real(Out22Real), 
    .Out22Imag(Out22Imag), 
    .Out23Real(Out23Real), 
    .Out23Imag(Out23Imag), 
    .Out24Real(Out24Real), 
    .Out24Imag(Out24Imag), 
    .Out31Real(Out31Real), 
    .Out31Imag(Out31Imag), 
    .Out32Real(Out32Real), 
    .Out32Imag(Out32Imag), 
    .Out33Real(Out33Real), 
    .Out33Imag(Out33Imag), 
    .Out34Real(Out34Real), 
    .Out34Imag(Out34Imag), 
    .Out41Real(Out41Real), 
    .Out41Imag(Out41Imag), 
    .Out42Real(Out42Real), 
    .Out42Imag(Out42Imag), 
    .Out43Real(Out43Real), 
    .Out43Imag(Out43Imag), 
    .Out44Real(Out44Real), 
    .Out44Imag(Out44Imag), 
    .OutMux(readdata)
    );



	// Instantiate the module
	RegistrodeListo RegistrodeListocopia (
    .CLK(clk),
    .ResetMaster(reset_n),
	 .Address(address),
    .EnableListo(EnableListo),
    .Out(OutInt),
    .Write(write)
    );





endmodule
