`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:02:04 12/01/2014 
// Design Name: 
// Module Name:    MainProyectoFinalPrueba 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MainProyectoFinal #(parameter Width = 32, ConLimitador=0,Magnitud = 7, Precision = 24, Signo = 1/*,
A00=  32'sb11110010000000000000000000000000, A01=  32'sb11110010100000000000000000000000, 
A02 =  32'sb11110011000000000000000000000000, A03 =  32'sb11110011100000000000000000000000, A04 =  32'sb11110100000000000000000000000000, A05 =  32'sb11110100100000000000000000000000, A06 =  32'sb11110101000000000000000000000000, A07 =  32'sb11110101100000000000000000000000, A08 =  32'sb11110110000000000000000000000000, A09 =  32'sb11110110100000000000000000000000,
A10=  32'sb11110111000000000000000000000000, A11=  32'sb11110111100000000000000000000000, A12 =  32'sb11111000000000000000000000000000, A13 =  32'sb11111000100000000000000000000000, A14 =  32'sb11111001000000000000000000000000, A15 =  32'sb11111001100000000000000000000000, A16 =  32'sb11111010000000000000000000000000, A17 =  32'sb11111010100000000000000000000000, A18 =  32'sb11111011000000000000000000000000, A19 =  32'sb11111011100000000000000000000000,
A20=  32'sb11111100000000000000000000000000, A21=  32'sb11111100100000000000000000000000, 
A22 =  32'sb11111101000000000000000000000000, A23 =  32'sb11111101100000000000000000000000, A24 =  32'sb11111110000000000000000000000000, A25 =  32'sb11111110100000000000000000000000, A26 =  32'sb11111111000000000000000000000000, A27 = 32'sb00000001000000000000000000000000, A28 = 32'sb00000011000000000000000000000000, A29 = 32'sb00001000000000000000000000000000, 
A30 = 32'sb00010100000000000000000000000000, 
M01= 32'sb00000000000000000000000000010010,  M02 = 32'sb00000000000000000000000000011101, M03 = 32'sb00000000000000000000000000110000, M04 = 32'sb00000000000000000000000001010000, M05 = 32'sb00000000000000000000000010000101, M06 = 32'sb00000000000000000000000011011011, M07 = 32'sb00000000000000000000000101101010, M08 = 32'sb00000000000000000000001001010100, M09 = 32'sb00000000000000000000001111011000, M10= 32'sb00000000000000000000011001010110, 
M11= 32'sb00000000000000000000101001110010, M12 = 32'sb00000000000000000001000100111000, M13 = 32'sb00000000000000000001110001100001, M14 = 32'sb00000000000000000010111011000100, M15 = 32'sb00000000000000000100110100001000, M16 = 32'sb00000000000000000111111011001110, M17 = 32'sb00000000000000001101000010001010, M18 = 32'sb00000000000000010101011001100010, M19 = 32'sb00000000000000100011000010100000, M20= 32'sb00000000000000111001000111101101, 
M21= 32'sb00000000000001011100011100110110,M22 = 32'sb00000000000010010011111001111110, M23 = 32'sb00000000000011101000010010000010, M24 = 32'sb00000000000101100010010111111111, M25 = 32'sb00000000001000000101011001111001, M26 = 32'sb00000000001011000100110111000010, M27 = 32'sb00000000001111010000001011111101, M28 = 32'sb00000000000110111100101101110000, M29 = 32'sb00000000000000011100111000110000,  M30 = 32'sb00000000000000000000000011000011,
B01= 32'sb00000000000000000000000100001001,  B02 = 32'sb00000000000000000000000110100111, B03 = 32'sb00000000000000000000001010100001, B04 = 32'sb00000000000000000000010000101110, B05 = 32'sb00000000000000000000011010100010, B06 = 32'sb00000000000000000000101010000010, B07 = 32'sb00000000000000000001000010011111, B08 = 32'sb00000000000000000001000010011111, B09 = 32'sb00000000000000000010100101010110,
B10= 32'sb00000000000000000100000011111011, B11= 32'sb00000000000000000110010111100110, B12 = 32'sb00000000000000001001111101011100, B13 = 32'sb00000000000000001111100001110111, B14 = 32'sb00000000000000011000001000001100, B15 = 32'sb00000000000000100101010101101000, B16 = 32'sb00000000000000111001100000100001, B17 = 32'sb00000000000001011000000100101101, B18 = 32'sb00000000000010000101111100100110, B19 = 32'sb00000000000011001001111011010011,
B20= 32'sb00000000000100101100111100011001, B21= 32'sb00000000000110111001101110001101,B22 = 32'sb00000000001001111011000000011110, B23 = 32'sb00000000001101110111000000110110, B24 = 32'sb00000000010010100110110111111101, B25 = 32'sb00000000010111101011101001001001, B26 = 32'sb00000000011100001010010101101101, B27 = 32'sb00000000100000000000000000000000, B28 = 32'sb00000000101001101000100000110000, B29 = 32'sb00000000111100111001100101111101, 
B30 = 32'sb00000000111111111111001101111011*/)
(CLK,MasterReset,write,read,address,writedata,readdata);
	 
	 
	 input CLK;
	 input MasterReset;
	 input write;	 
	 input read;
	 input [8:0] address;
	 input signed [Width-1:0] writedata;
	 output signed [Width-1:0] readdata;
	 
	 wire ResetInterfaz,ResetStart,ResetCoeffALUandInput,       
	  EnableCoeffALUandInput,EnableMulX,EnableRegOutMultCoeffX,EnableFuctAct,EnableRegActFunc,
	  EnableMulY,EnableRegDesplazamiento,EnableSum,SELOffset,EnableAcumulador,ResetAcumulador,
	  Listo,Start,Error1;
	  
	  wire signed [Width-1:0] Coeff00,Coeff01,Coeff02,Coeff03,Coeff04,Coeff05,Coeff06,Coeff07,Coeff08,
	  Coeff09,Coeff10,Coeff11,Coeff12,Coeff13,Coeff14,Coeff15,Coeff16,Coeff17,Coeff18,Coeff19,Offset,
	  InDato,InDatoALU,Acumulador,OutALU,Y0,Y1,Y2,Y3,Y4,Y5,Y6,Y7,Y8,Y9;
	  
	  wire [3:0] SELCoeffY,SELCoeffX;
	  
	  reg Error;
	 
	 FSMNeuralNetwork FSMNeuralNetworkCopia (
    .CLK(CLK),                        //**********************************
    .reset(~MasterReset),              //**********************************
    .Start(Start),                    //**********************************
    .Read(read),                      //**********************************
    .Address(address),                //**********************************
    .ResetInterfaz(ResetInterfaz),    //**********************************
    .ResetStart(ResetStart),          //**********************************
    .ResetCoeffALUandInput(ResetCoeffALUandInput),  //**********************************
    .EnableCoeffALUandInput(EnableCoeffALUandInput),    //**********************************
    .EnableMulX(EnableMulX),                           //**********************************
    .SELCoeffX(SELCoeffX),                             //**********************************
    .EnableRegOutMultCoeffX(EnableRegOutMultCoeffX),      //********************************** 
    .EnableFuctAct(EnableFuctAct),                      //**********************************
    .EnableRegActFunc(EnableRegActFunc),                 //**********************************
    .EnableMulY(EnableMulY),                              //**********************************
    .EnableRegDesplazamiento(EnableRegDesplazamiento),    //**********************************
    .EnableSum(EnableSum),                               //**********************************
    .SELCoeffY(SELCoeffY),                              //**********************************
    .SELOffset(SELOffset),                              //**********************************
    .EnableAcumulador(EnableAcumulador),                //**********************************
    .ResetAcumulador(ResetAcumulador),                   //**********************************
    .Listo(Listo)                                       //**********************************
    );
	 
	 
	 
	 
	 RegistroCargaInterfaz   #(.Width(Width)) RegistroCargaInterfazCopia (
    .CLK(CLK),                               //**********************************
    .Reset(ResetInterfaz),                   //**********************************
    .ResetStart(ResetStart),                 //**********************************
    .InDatoMemoria(writedata),               //********************************** 
    .Write(write),                           //********************************** 
    .Address(address),                       //********************************** 
    .Coeff00(Coeff00),                       //**********************************
    .Coeff01(Coeff01),                       //**********************************
    .Coeff02(Coeff02),                       //**********************************
    .Coeff03(Coeff03),                       //**********************************
    .Coeff04(Coeff04),                       //**********************************
    .Coeff05(Coeff05),                       //**********************************
    .Coeff06(Coeff06),                       //**********************************
    .Coeff07(Coeff07),                       //********************************** 
    .Coeff08(Coeff08),                       //**********************************
    .Coeff09(Coeff09),                       //********************************** 
    .Coeff10(Coeff10),                       //**********************************
    .Coeff11(Coeff11),                       //**********************************
    .Coeff12(Coeff12),                       //********************************** 
    .Coeff13(Coeff13),                       //********************************** 
    .Coeff14(Coeff14),                       //********************************** 
    .Coeff15(Coeff15),                       //**********************************
    .Coeff16(Coeff16),                       //**********************************
    .Coeff17(Coeff17),                       //********************************** 
    .Coeff18(Coeff18),                       //**********************************
    .Coeff19(Coeff19),                       //**********************************
    .Offset(Offset),                         //**********************************
    .InDato(InDato),                         //**********************************
    .Start(Start)                            //**********************************
    );
	 
	 Registro  #(.Width(Width)) RegistroEntrada (
    .CLK(CLK),                               //**********************************
    .reset(ResetCoeffALUandInput),           //**********************************
    .Enable(EnableCoeffALUandInput),         //**********************************
    .Entrada(InDato),                        //**********************************
    .Salida(InDatoALU)                       //**********************************
    );
	 
	 ALUNeuralNetwork #(.Width(Width),.Magnitud(Magnitud),.ConLimitador(ConLimitador),.Precision(Precision), .Signo(Signo), 
	   /*.A00(A00), 
		.A01(A01),.A02(A02),.A03(A03),.A04(A04),.A05(A05),.A06(A06),.A07(A07),.A08(A08),.A09(A09),
		.A10(A10),.A11(A11),.A12(A12),.A13(A13),.A14(A14),.A15(A15),.A16(A16),.A17(A17),.A18(A18),.A19(A19),
		.A20(A20),.A21(A21),.A22(A22),.A23(A23),.A24(A24),.A25(A25),.A26(A26),.A27(A27),.A28(A28),.A29(A29), 
		.A30(A30), 
		.M01(M01),.M02(M02),.M03(M03),.M04(M04),.M05(M05),.M06(M06),.M07(M07),.M08(M08),.M09(M09),
		.M10(M10),.M11(M11),.M12(M12),.M13(M13),.M14(M14),.M15(M15),.M16(M16),.M17(M17),.M18(M18),.M19(M19),
		.M20(M20),.M21(M21),.M22(M22),.M23(M23),.M24(M24),.M25(M25),.M26(M26),.M27(M27),.M28(M28),.M29(M29), 
		.M30(M30),
		.B01(B01),.B02(B02),.B03(B03),.B04(B04),.B05(B05),.B06(B06),.B07(B07),.B08(B08),.B09(B09),
		.B10(B10),.B11(B11),.B12(B12),.B13(B13),.B14(B14),.B15(B15),.B16(B16),.B17(B17),.B18(B18),.B19(B19),
		.B20(B20),.B21(B21),.B22(B22),.B23(B23),.B24(B24),.B25(B25),.B26(B26),.B27(B27),.B28(B28),.B29(B29), 
		.B30(B30)*/
		.A00(32'sb11110010000000000000000000000000), .A01(32'sb11110010100000000000000000000000), 
		.A02(32'sb11110011000000000000000000000000), .A03(32'sb11110011100000000000000000000000), .A04(32'sb11110100000000000000000000000000), .A05(32'sb11110100100000000000000000000000), .A06(32'sb11110101000000000000000000000000), .A07(32'sb11110101100000000000000000000000), .A08(32'sb11110110000000000000000000000000), .A09(32'sb11110110100000000000000000000000),
		.A10(32'sb11110111000000000000000000000000), .A11(32'sb11110111100000000000000000000000), .A12(32'sb11111000000000000000000000000000), .A13(32'sb11111000100000000000000000000000), .A14(32'sb11111001000000000000000000000000), .A15(32'sb11111001100000000000000000000000), .A16(32'sb11111010000000000000000000000000), .A17(32'sb11111010100000000000000000000000), .A18(32'sb11111011000000000000000000000000), .A19(32'sb11111011100000000000000000000000),
		.A20(32'sb11111100000000000000000000000000), .A21(32'sb11111100100000000000000000000000), 
		.A22(32'sb11111101000000000000000000000000), .A23(32'sb11111101100000000000000000000000), .A24(32'sb11111110000000000000000000000000), .A25(32'sb11111110100000000000000000000000), .A26(32'sb11111111000000000000000000000000), .A27(32'sb00000001000000000000000000000000), .A28(32'sb00000011000000000000000000000000), .A29(32'sb00001000000000000000000000000000), 
		.A30(32'sb00010100000000000000000000000000), 
		.M01(32'sb00000000000000000000000000010010), .M02(32'sb00000000000000000000000000011101), .M03(32'sb00000000000000000000000000110000), .M04(32'sb00000000000000000000000001010000), .M05(32'sb00000000000000000000000010000101), .M06(32'sb00000000000000000000000011011011), .M07(32'sb00000000000000000000000101101010), .M08(32'sb00000000000000000000001001010100), .M09(32'sb00000000000000000000001111011000), .M10(32'sb00000000000000000000011001010110), 
		.M11(32'sb00000000000000000000101001110010), .M12(32'sb00000000000000000001000100111000), .M13(32'sb00000000000000000001110001100001), .M14(32'sb00000000000000000010111011000100), .M15(32'sb00000000000000000100110100001000), .M16(32'sb00000000000000000111111011001110), .M17(32'sb00000000000000001101000010001010), .M18(32'sb00000000000000010101011001100010), .M19(32'sb00000000000000100011000010100000), .M20(32'sb00000000000000111001000111101101), 
		.M21(32'sb00000000000001011100011100110110), .M22(32'sb00000000000010010011111001111110), .M23(32'sb00000000000011101000010010000010), .M24(32'sb00000000000101100010010111111111), .M25(32'sb00000000001000000101011001111001), .M26(32'sb00000000001011000100110111000010), .M27(32'sb00000000001111010000001011111101), .M28(32'sb00000000000110111100101101110000), .M29(32'sb00000000000000011100111000110000), .M30(32'sb00000000000000000000000011000011),
		.B01(32'sb00000000000000000000000100001001), .B02(32'sb00000000000000000000000110100111), .B03(32'sb00000000000000000000001010100001), .B04(32'sb00000000000000000000010000101110), .B05(32'sb00000000000000000000011010100010), .B06(32'sb00000000000000000000101010000010), .B07(32'sb00000000000000000001000010011111), .B08(32'sb00000000000000000001000010011111), .B09(32'sb00000000000000000010100101010110),
		.B10(32'sb00000000000000000100000011111011), .B11(32'sb00000000000000000110010111100110), .B12(32'sb00000000000000001001111101011100), .B13(32'sb00000000000000001111100001110111), .B14(32'sb00000000000000011000001000001100), .B15(32'sb00000000000000100101010101101000), .B16(32'sb00000000000000111001100000100001), .B17(32'sb00000000000001011000000100101101), .B18(32'sb00000000000010000101111100100110), .B19(32'sb00000000000011001001111011010011),
		.B20(32'sb00000000000100101100111100011001), .B21(32'sb00000000000110111001101110001101), .B22(32'sb00000000001001111011000000011110), .B23(32'sb00000000001101110111000000110110), .B24(32'sb00000000010010100110110111111101), .B25(32'sb00000000010111101011101001001001), .B26(32'sb00000000011100001010010101101101), .B27(32'sb00000000100000000000000000000000), .B28(32'sb00000000101001101000100000110000), .B29(32'sb00000000111100111001100101111101), 
		.B30(32'sb00000000111111111111001101111011)
		)
	 ALUNeuralNetworkCopia (
    .CLK(CLK),                                //**********************************
    .reset(ResetCoeffALUandInput),             //**********************************
    .EnableLoadCoeff(EnableCoeffALUandInput),         //**********************************
    .EnableMulX(EnableMulX),                   //**********************************
    .EnableRegOutMultCoeffX(EnableRegOutMultCoeffX), //**********************************
    .EnableFuctAct(EnableFuctAct),                   //**********************************
    .EnableRegActFunc(EnableRegActFunc),             //********************************** 
    .EnableMulY(EnableMulY),                          //**********************************
    .EnableRegDesplazamiento(EnableRegDesplazamiento),    //**********************************
    .EnableSum(EnableSum),                                  //**********************************
    .InDato(InDatoALU),                       //**********************************
    .Acumulador(Acumulador),                  //**********************************
    .SELCoeffX(SELCoeffX),                     //**********************************
    .SELCoeffY(SELCoeffY),                     //**********************************
    .SELOffset(SELOffset),                    //**********************************
    .Coeff00(Coeff00),                        //**********************************
    .Coeff01(Coeff01),                        //**********************************
    .Coeff02(Coeff02),                        //**********************************
    .Coeff03(Coeff03),                        //**********************************
    .Coeff04(Coeff04),                        //**********************************
    .Coeff05(Coeff05),                        //**********************************
    .Coeff06(Coeff06),                        //**********************************
    .Coeff07(Coeff07),                         //**********************************
    .Coeff08(Coeff08),                        //********************************** 
    .Coeff09(Coeff09),                        //********************************** 
    .Coeff10(Coeff10),                         //********************************** 
    .Coeff11(Coeff11),                        //**********************************
    .Coeff12(Coeff12),                        //**********************************
    .Coeff13(Coeff13),                           //**********************************
    .Coeff14(Coeff14),                           //**********************************
    .Coeff15(Coeff15),                          //**********************************
    .Coeff16(Coeff16),                           //**********************************
    .Coeff17(Coeff17),                          //**********************************
    .Coeff18(Coeff18),                          //**********************************
    .Coeff19(Coeff19),                            //**********************************
    .Offset(Offset),                            //**********************************
    .Error(Error1),                             //**********************************
    .OutDato(OutALU),                           //**********************************
    .Y0(Y0),                                    //**********************************
    .Y1(Y1),                                    //**********************************
    .Y2(Y2),                                    //**********************************
    .Y3(Y3),                                    //**********************************
    .Y4(Y4),                                    //**********************************
    .Y5(Y5),                                    //**********************************
    .Y6(Y6),                                    //**********************************
    .Y7(Y7),                                    //**********************************
    .Y8(Y8),                                    //**********************************
    .Y9(Y9)                                     //**********************************
    );
	 
	 Registro  #(.Width(Width)) RegistroAcumulador (
    .CLK(CLK),                           //**********************************
    .reset(ResetAcumulador),             //**********************************
    .Enable(EnableAcumulador),           //**********************************
    .Entrada(OutALU),                    //**********************************
    .Salida(Acumulador)                  //**********************************
    );
	 
	 EscrituraRegistroToMemoria  #(.Width(Width)) EscrituraRegistroToMemoriaPruebaCopia (
    .Read(read),                     //**********************************
    .InError(Error),                 //**********************************
    .Address(address),               //**********************************
    .ListoIn(Listo),                 //**********************************
    .InDato(Acumulador),             //**********************************
    .Coeff00(Coeff00),               //**********************************
    .Coeff01(Coeff01),               //**********************************
    .Coeff02(Coeff02),               //**********************************
    .Coeff03(Coeff03),               //**********************************
    .Coeff04(Coeff04),               //********************************** 
    .Coeff05(Coeff05),               //********************************** 
    .Coeff06(Coeff06),               //********************************** 
    .Coeff07(Coeff07),               //********************************** 
    .Coeff08(Coeff08),               //********************************** 
    .Coeff09(Coeff09),               //********************************** 
    .Coeff10(Coeff10),               //**********************************
    .Coeff11(Coeff11),               //**********************************
    .Coeff12(Coeff12),               //**********************************
    .Coeff13(Coeff13),               //**********************************
    .Coeff14(Coeff14),               //********************************** 
    .Coeff15(Coeff15),               //********************************** 
    .Coeff16(Coeff16),               //********************************** 
    .Coeff17(Coeff17),               //**********************************
    .Coeff18(Coeff18),               //**********************************
    .Coeff19(Coeff19),               //**********************************
    .Offset(Offset),                 //**********************************
    .DatoEntradaSistema(InDatoALU),  //**********************************
    .Y0(Y0),                         //**********************************
    .Y1(Y1),                          //**********************************
    .Y2(Y2),                         //**********************************
    .Y3(Y3),                         //**********************************
    .Y4(Y4),                         //********************************** 
    .Y5(Y5),                         //**********************************
    .Y6(Y6),                         //**********************************
    .Y7(Y7),                         //**********************************
    .Y8(Y8),                         //**********************************
    .Y9(Y9),                         //**********************************
    .OutDato(readdata)              //**********************************
    );
	 
	 
	 always @(posedge CLK) begin  //***************REGISTRO QUE ALMACENA EN CASO DE QUE HAYA ERRORES
      if (ResetStart) begin
         Error <= 1'b0;
      end else if (Error1) begin
         Error <= 1'b1;
      end
	 end





endmodule
