// SOC.v

// Generated using ACDS version 13.0sp1 232 at 2014.11.27.23:14:43

`timescale 1 ps / 1 ps
module SOC (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         nios_ii_instruction_master_waitrequest;                                                             // NIOS_II_instruction_master_translator:av_waitrequest -> NIOS_II:i_waitrequest
	wire  [15:0] nios_ii_instruction_master_address;                                                                 // NIOS_II:i_address -> NIOS_II_instruction_master_translator:av_address
	wire         nios_ii_instruction_master_read;                                                                    // NIOS_II:i_read -> NIOS_II_instruction_master_translator:av_read
	wire  [31:0] nios_ii_instruction_master_readdata;                                                                // NIOS_II_instruction_master_translator:av_readdata -> NIOS_II:i_readdata
	wire         nios_ii_data_master_waitrequest;                                                                    // NIOS_II_data_master_translator:av_waitrequest -> NIOS_II:d_waitrequest
	wire  [31:0] nios_ii_data_master_writedata;                                                                      // NIOS_II:d_writedata -> NIOS_II_data_master_translator:av_writedata
	wire  [15:0] nios_ii_data_master_address;                                                                        // NIOS_II:d_address -> NIOS_II_data_master_translator:av_address
	wire         nios_ii_data_master_write;                                                                          // NIOS_II:d_write -> NIOS_II_data_master_translator:av_write
	wire         nios_ii_data_master_read;                                                                           // NIOS_II:d_read -> NIOS_II_data_master_translator:av_read
	wire  [31:0] nios_ii_data_master_readdata;                                                                       // NIOS_II_data_master_translator:av_readdata -> NIOS_II:d_readdata
	wire         nios_ii_data_master_debugaccess;                                                                    // NIOS_II:jtag_debug_module_debugaccess_to_roms -> NIOS_II_data_master_translator:av_debugaccess
	wire   [3:0] nios_ii_data_master_byteenable;                                                                     // NIOS_II:d_byteenable -> NIOS_II_data_master_translator:av_byteenable
	wire         nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                               // NIOS_II:jtag_debug_module_waitrequest -> NIOS_II_jtag_debug_module_translator:av_waitrequest
	wire  [31:0] nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                 // NIOS_II_jtag_debug_module_translator:av_writedata -> NIOS_II:jtag_debug_module_writedata
	wire   [8:0] nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_address;                                   // NIOS_II_jtag_debug_module_translator:av_address -> NIOS_II:jtag_debug_module_address
	wire         nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_write;                                     // NIOS_II_jtag_debug_module_translator:av_write -> NIOS_II:jtag_debug_module_write
	wire         nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_read;                                      // NIOS_II_jtag_debug_module_translator:av_read -> NIOS_II:jtag_debug_module_read
	wire  [31:0] nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                  // NIOS_II:jtag_debug_module_readdata -> NIOS_II_jtag_debug_module_translator:av_readdata
	wire         nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                               // NIOS_II_jtag_debug_module_translator:av_debugaccess -> NIOS_II:jtag_debug_module_debugaccess
	wire   [3:0] nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                // NIOS_II_jtag_debug_module_translator:av_byteenable -> NIOS_II:jtag_debug_module_byteenable
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_writedata;                                                    // RAM_s1_translator:av_writedata -> RAM:writedata
	wire  [11:0] ram_s1_translator_avalon_anti_slave_0_address;                                                      // RAM_s1_translator:av_address -> RAM:address
	wire         ram_s1_translator_avalon_anti_slave_0_chipselect;                                                   // RAM_s1_translator:av_chipselect -> RAM:chipselect
	wire         ram_s1_translator_avalon_anti_slave_0_clken;                                                        // RAM_s1_translator:av_clken -> RAM:clken
	wire         ram_s1_translator_avalon_anti_slave_0_write;                                                        // RAM_s1_translator:av_write -> RAM:write
	wire  [31:0] ram_s1_translator_avalon_anti_slave_0_readdata;                                                     // RAM:readdata -> RAM_s1_translator:av_readdata
	wire   [3:0] ram_s1_translator_avalon_anti_slave_0_byteenable;                                                   // RAM_s1_translator:av_byteenable -> RAM:byteenable
	wire         ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                          // Ifsr_0_avalon_slave_0_translator:av_read -> Ifsr_0:read
	wire  [31:0] ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                                      // Ifsr_0:read_data -> Ifsr_0_avalon_slave_0_translator:av_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                           // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                             // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                               // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                            // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                 // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                              // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [0:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                  // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                 // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                  // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                               // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                    // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                 // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_waitrequest;                        // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_II_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios_ii_instruction_master_translator_avalon_universal_master_0_burstcount;                         // NIOS_II_instruction_master_translator:uav_burstcount -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios_ii_instruction_master_translator_avalon_universal_master_0_writedata;                          // NIOS_II_instruction_master_translator:uav_writedata -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [15:0] nios_ii_instruction_master_translator_avalon_universal_master_0_address;                            // NIOS_II_instruction_master_translator:uav_address -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_lock;                               // NIOS_II_instruction_master_translator:uav_lock -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_write;                              // NIOS_II_instruction_master_translator:uav_write -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_read;                               // NIOS_II_instruction_master_translator:uav_read -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios_ii_instruction_master_translator_avalon_universal_master_0_readdata;                           // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_II_instruction_master_translator:uav_readdata
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_debugaccess;                        // NIOS_II_instruction_master_translator:uav_debugaccess -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios_ii_instruction_master_translator_avalon_universal_master_0_byteenable;                         // NIOS_II_instruction_master_translator:uav_byteenable -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_readdatavalid;                      // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_II_instruction_master_translator:uav_readdatavalid
	wire         nios_ii_data_master_translator_avalon_universal_master_0_waitrequest;                               // NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> NIOS_II_data_master_translator:uav_waitrequest
	wire   [2:0] nios_ii_data_master_translator_avalon_universal_master_0_burstcount;                                // NIOS_II_data_master_translator:uav_burstcount -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios_ii_data_master_translator_avalon_universal_master_0_writedata;                                 // NIOS_II_data_master_translator:uav_writedata -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [15:0] nios_ii_data_master_translator_avalon_universal_master_0_address;                                   // NIOS_II_data_master_translator:uav_address -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios_ii_data_master_translator_avalon_universal_master_0_lock;                                      // NIOS_II_data_master_translator:uav_lock -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios_ii_data_master_translator_avalon_universal_master_0_write;                                     // NIOS_II_data_master_translator:uav_write -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios_ii_data_master_translator_avalon_universal_master_0_read;                                      // NIOS_II_data_master_translator:uav_read -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios_ii_data_master_translator_avalon_universal_master_0_readdata;                                  // NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_readdata -> NIOS_II_data_master_translator:uav_readdata
	wire         nios_ii_data_master_translator_avalon_universal_master_0_debugaccess;                               // NIOS_II_data_master_translator:uav_debugaccess -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios_ii_data_master_translator_avalon_universal_master_0_byteenable;                                // NIOS_II_data_master_translator:uav_byteenable -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios_ii_data_master_translator_avalon_universal_master_0_readdatavalid;                             // NIOS_II_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> NIOS_II_data_master_translator:uav_readdatavalid
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // NIOS_II_jtag_debug_module_translator:uav_waitrequest -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> NIOS_II_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                   // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> NIOS_II_jtag_debug_module_translator:uav_writedata
	wire  [15:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                     // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> NIOS_II_jtag_debug_module_translator:uav_address
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                       // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> NIOS_II_jtag_debug_module_translator:uav_write
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                        // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> NIOS_II_jtag_debug_module_translator:uav_lock
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                        // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> NIOS_II_jtag_debug_module_translator:uav_read
	wire  [31:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                    // NIOS_II_jtag_debug_module_translator:uav_readdata -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // NIOS_II_jtag_debug_module_translator:uav_readdatavalid -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> NIOS_II_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> NIOS_II_jtag_debug_module_translator:uav_byteenable
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                 // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // RAM_s1_translator:uav_waitrequest -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // RAM_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> RAM_s1_translator:uav_burstcount
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // RAM_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> RAM_s1_translator:uav_writedata
	wire  [15:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // RAM_s1_translator_avalon_universal_slave_0_agent:m0_address -> RAM_s1_translator:uav_address
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // RAM_s1_translator_avalon_universal_slave_0_agent:m0_write -> RAM_s1_translator:uav_write
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // RAM_s1_translator_avalon_universal_slave_0_agent:m0_lock -> RAM_s1_translator:uav_lock
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // RAM_s1_translator_avalon_universal_slave_0_agent:m0_read -> RAM_s1_translator:uav_read
	wire  [31:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // RAM_s1_translator:uav_readdata -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // RAM_s1_translator:uav_readdatavalid -> RAM_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> RAM_s1_translator:uav_debugaccess
	wire   [3:0] ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // RAM_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> RAM_s1_translator:uav_byteenable
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // RAM_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // Ifsr_0_avalon_slave_0_translator:uav_waitrequest -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Ifsr_0_avalon_slave_0_translator:uav_burstcount
	wire  [31:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Ifsr_0_avalon_slave_0_translator:uav_writedata
	wire  [15:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                         // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Ifsr_0_avalon_slave_0_translator:uav_address
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                           // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Ifsr_0_avalon_slave_0_translator:uav_write
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                            // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Ifsr_0_avalon_slave_0_translator:uav_lock
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                            // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Ifsr_0_avalon_slave_0_translator:uav_read
	wire  [31:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // Ifsr_0_avalon_slave_0_translator:uav_readdata -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // Ifsr_0_avalon_slave_0_translator:uav_readdatavalid -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Ifsr_0_avalon_slave_0_translator:uav_debugaccess
	wire   [3:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Ifsr_0_avalon_slave_0_translator:uav_byteenable
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [15:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire  [15:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [15:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [89:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [89:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                     // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [88:0] nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                      // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router:sink_ready -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // NIOS_II_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_valid;                            // NIOS_II_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // NIOS_II_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [88:0] nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_data;                             // NIOS_II_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_001:sink_ready -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                       // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [88:0] nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                        // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router:sink_ready -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // RAM_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // RAM_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // RAM_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [88:0] ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // RAM_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_001:sink_ready -> RAM_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                           // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [88:0] ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                            // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [88:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [88:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_004:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [88:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_005:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                                     // rst_controller:reset_out -> [Ifsr_0:rst_n, Ifsr_0_avalon_slave_0_translator:reset, Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, NIOS_II:reset_n, NIOS_II_data_master_translator:reset, NIOS_II_data_master_translator_avalon_universal_master_0_agent:reset, NIOS_II_instruction_master_translator:reset, NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:reset, NIOS_II_jtag_debug_module_translator:reset, NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, RAM:reset, RAM_s1_translator:reset, RAM_s1_translator_avalon_universal_slave_0_agent:reset, RAM_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         rst_controller_reset_out_reset_req;                                                                 // rst_controller:reset_req -> RAM:reset_req
	wire         cmd_xbar_demux_src0_endofpacket;                                                                    // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                          // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                  // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src0_data;                                                                           // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [5:0] cmd_xbar_demux_src0_channel;                                                                        // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                          // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                    // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                          // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                  // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src1_data;                                                                           // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [5:0] cmd_xbar_demux_src1_channel;                                                                        // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                          // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_src2_endofpacket;                                                                    // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                          // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                  // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [88:0] cmd_xbar_demux_src2_data;                                                                           // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [5:0] cmd_xbar_demux_src2_channel;                                                                        // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire         cmd_xbar_demux_src2_ready;                                                                          // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                      // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                              // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src0_data;                                                                       // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src0_channel;                                                                    // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                      // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                      // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                              // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src1_data;                                                                       // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src1_channel;                                                                    // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                      // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                      // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                              // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src2_data;                                                                       // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src2_channel;                                                                    // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire         cmd_xbar_demux_001_src2_ready;                                                                      // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                                // cmd_xbar_demux_001:src3_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                      // cmd_xbar_demux_001:src3_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                              // cmd_xbar_demux_001:src3_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src3_data;                                                                       // cmd_xbar_demux_001:src3_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src3_channel;                                                                    // cmd_xbar_demux_001:src3_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                                // cmd_xbar_demux_001:src4_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                      // cmd_xbar_demux_001:src4_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                              // cmd_xbar_demux_001:src4_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src4_data;                                                                       // cmd_xbar_demux_001:src4_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src4_channel;                                                                    // cmd_xbar_demux_001:src4_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                                // cmd_xbar_demux_001:src5_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                      // cmd_xbar_demux_001:src5_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                              // cmd_xbar_demux_001:src5_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_demux_001_src5_data;                                                                       // cmd_xbar_demux_001:src5_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src5_channel;                                                                    // cmd_xbar_demux_001:src5_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                    // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                          // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                  // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [88:0] rsp_xbar_demux_src0_data;                                                                           // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [5:0] rsp_xbar_demux_src0_channel;                                                                        // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                          // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                    // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                          // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                  // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [88:0] rsp_xbar_demux_src1_data;                                                                           // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [5:0] rsp_xbar_demux_src1_channel;                                                                        // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                          // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                      // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                              // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src0_data;                                                                       // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src0_channel;                                                                    // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                      // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                      // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                              // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [88:0] rsp_xbar_demux_001_src1_data;                                                                       // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src1_channel;                                                                    // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                      // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                      // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                              // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [88:0] rsp_xbar_demux_002_src0_data;                                                                       // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [5:0] rsp_xbar_demux_002_src0_channel;                                                                    // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                      // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_002_src1_endofpacket;                                                                // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src1_valid;                                                                      // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src1_startofpacket;                                                              // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [88:0] rsp_xbar_demux_002_src1_data;                                                                       // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [5:0] rsp_xbar_demux_002_src1_channel;                                                                    // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src1_ready;                                                                      // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                      // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                              // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [88:0] rsp_xbar_demux_003_src0_data;                                                                       // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire   [5:0] rsp_xbar_demux_003_src0_channel;                                                                    // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                      // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                      // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                              // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [88:0] rsp_xbar_demux_004_src0_data;                                                                       // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [5:0] rsp_xbar_demux_004_src0_channel;                                                                    // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                      // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                      // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                              // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [88:0] rsp_xbar_demux_005_src0_data;                                                                       // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [5:0] rsp_xbar_demux_005_src0_channel;                                                                    // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                      // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         addr_router_src_endofpacket;                                                                        // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                              // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                      // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [88:0] addr_router_src_data;                                                                               // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [5:0] addr_router_src_channel;                                                                            // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                              // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                       // rsp_xbar_mux:src_endofpacket -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                             // rsp_xbar_mux:src_valid -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                     // rsp_xbar_mux:src_startofpacket -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] rsp_xbar_mux_src_data;                                                                              // rsp_xbar_mux:src_data -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] rsp_xbar_mux_src_channel;                                                                           // rsp_xbar_mux:src_channel -> NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                             // NIOS_II_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                    // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                          // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                  // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [88:0] addr_router_001_src_data;                                                                           // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [5:0] addr_router_001_src_channel;                                                                        // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                          // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                   // rsp_xbar_mux_001:src_endofpacket -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                         // rsp_xbar_mux_001:src_valid -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                 // rsp_xbar_mux_001:src_startofpacket -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [88:0] rsp_xbar_mux_001_src_data;                                                                          // rsp_xbar_mux_001:src_data -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] rsp_xbar_mux_001_src_channel;                                                                       // rsp_xbar_mux_001:src_channel -> NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                         // NIOS_II_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                       // cmd_xbar_mux:src_endofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                             // cmd_xbar_mux:src_valid -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                     // cmd_xbar_mux:src_startofpacket -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_src_data;                                                                              // cmd_xbar_mux:src_data -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_src_channel;                                                                           // cmd_xbar_mux:src_channel -> NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                             // NIOS_II_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                          // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                        // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [88:0] id_router_src_data;                                                                                 // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [5:0] id_router_src_channel;                                                                              // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                   // cmd_xbar_mux_001:src_endofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                         // cmd_xbar_mux_001:src_valid -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                 // cmd_xbar_mux_001:src_startofpacket -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_001_src_data;                                                                          // cmd_xbar_mux_001:src_data -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_001_src_channel;                                                                       // cmd_xbar_mux_001:src_channel -> RAM_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                         // RAM_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                      // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                            // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                    // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [88:0] id_router_001_src_data;                                                                             // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [5:0] id_router_001_src_channel;                                                                          // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                            // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_mux_002_src_endofpacket;                                                                   // cmd_xbar_mux_002:src_endofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_002_src_valid;                                                                         // cmd_xbar_mux_002:src_valid -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_002_src_startofpacket;                                                                 // cmd_xbar_mux_002:src_startofpacket -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [88:0] cmd_xbar_mux_002_src_data;                                                                          // cmd_xbar_mux_002:src_data -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_002_src_channel;                                                                       // cmd_xbar_mux_002:src_channel -> Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_002_src_ready;                                                                         // Ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire         id_router_002_src_endofpacket;                                                                      // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                            // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                    // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [88:0] id_router_002_src_data;                                                                             // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [5:0] id_router_002_src_channel;                                                                          // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                            // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                      // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                            // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                    // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [88:0] id_router_003_src_data;                                                                             // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [5:0] id_router_003_src_channel;                                                                          // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                            // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                      // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                      // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                            // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                    // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [88:0] id_router_004_src_data;                                                                             // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [5:0] id_router_004_src_channel;                                                                          // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                            // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                      // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                            // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                    // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [88:0] id_router_005_src_data;                                                                             // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [5:0] id_router_005_src_channel;                                                                          // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                            // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         irq_mapper_receiver0_irq;                                                                           // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                           // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_ii_d_irq_irq;                                                                                  // irq_mapper:sender_irq -> NIOS_II:d_irq

	SOC_RAM ram (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	SOC_NIOS_II nios_ii (
		.clk                                   (clk_clk),                                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                      //                   reset_n.reset_n
		.d_address                             (nios_ii_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios_ii_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios_ii_data_master_read),                                             //                          .read
		.d_readdata                            (nios_ii_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios_ii_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios_ii_data_master_write),                                            //                          .write
		.d_writedata                           (nios_ii_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_ii_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios_ii_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios_ii_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios_ii_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios_ii_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios_ii_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                     //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                      // custom_instruction_master.readra
	);

	SOC_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	SOC_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                                            //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                    //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	SOC_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                              //   irq.irq
	);

	lfsr ifsr_0 (
		.clk       (clk_clk),                                                       //          clock.clk
		.read      (ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read),     // avalon_slave_0.read
		.read_data (ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata), //               .readdata
		.rst_n     (~rst_controller_reset_out_reset)                                //   reset_sink_1.reset_n
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios_ii_instruction_master_translator (
		.clk                      (clk_clk),                                                                       //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                     reset.reset
		.uav_address              (nios_ii_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_ii_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_ii_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_ii_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_ii_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_ii_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_ii_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_ii_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_ii_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_ii_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_ii_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_ii_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_ii_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios_ii_instruction_master_read),                                               //                          .read
		.av_readdata              (nios_ii_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                          //               (terminated)
		.av_byteenable            (4'b1111),                                                                       //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                          //               (terminated)
		.av_begintransfer         (1'b0),                                                                          //               (terminated)
		.av_chipselect            (1'b0),                                                                          //               (terminated)
		.av_readdatavalid         (),                                                                              //               (terminated)
		.av_write                 (1'b0),                                                                          //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                          //               (terminated)
		.av_lock                  (1'b0),                                                                          //               (terminated)
		.av_debugaccess           (1'b0),                                                                          //               (terminated)
		.uav_clken                (),                                                                              //               (terminated)
		.av_clken                 (1'b1),                                                                          //               (terminated)
		.uav_response             (2'b00),                                                                         //               (terminated)
		.av_response              (),                                                                              //               (terminated)
		.uav_writeresponserequest (),                                                                              //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                          //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                          //               (terminated)
		.av_writeresponsevalid    ()                                                                               //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (16),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (16),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios_ii_data_master_translator (
		.clk                      (clk_clk),                                                                //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                     reset.reset
		.uav_address              (nios_ii_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios_ii_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios_ii_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios_ii_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios_ii_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios_ii_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios_ii_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios_ii_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios_ii_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios_ii_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios_ii_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios_ii_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios_ii_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios_ii_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios_ii_data_master_read),                                               //                          .read
		.av_readdata              (nios_ii_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios_ii_data_master_write),                                              //                          .write
		.av_writedata             (nios_ii_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios_ii_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                   //               (terminated)
		.av_begintransfer         (1'b0),                                                                   //               (terminated)
		.av_chipselect            (1'b0),                                                                   //               (terminated)
		.av_readdatavalid         (),                                                                       //               (terminated)
		.av_lock                  (1'b0),                                                                   //               (terminated)
		.uav_clken                (),                                                                       //               (terminated)
		.av_clken                 (1'b1),                                                                   //               (terminated)
		.uav_response             (2'b00),                                                                  //               (terminated)
		.av_response              (),                                                                       //               (terminated)
		.uav_writeresponserequest (),                                                                       //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                   //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                   //               (terminated)
		.av_writeresponsevalid    ()                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios_ii_jtag_debug_module_translator (
		.clk                      (clk_clk),                                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios_ii_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_chipselect            (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ram_s1_translator (
		.clk                      (clk_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //                    reset.reset
		.uav_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                  //              (terminated)
		.av_begintransfer         (),                                                                  //              (terminated)
		.av_beginbursttransfer    (),                                                                  //              (terminated)
		.av_burstcount            (),                                                                  //              (terminated)
		.av_readdatavalid         (1'b0),                                                              //              (terminated)
		.av_waitrequest           (1'b0),                                                              //              (terminated)
		.av_writebyteenable       (),                                                                  //              (terminated)
		.av_lock                  (),                                                                  //              (terminated)
		.uav_clken                (1'b0),                                                              //              (terminated)
		.av_debugaccess           (),                                                                  //              (terminated)
		.av_outputenable          (),                                                                  //              (terminated)
		.uav_response             (),                                                                  //              (terminated)
		.av_response              (2'b00),                                                             //              (terminated)
		.uav_writeresponserequest (1'b0),                                                              //              (terminated)
		.uav_writeresponsevalid   (),                                                                  //              (terminated)
		.av_writeresponserequest  (),                                                                  //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ifsr_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_read                  (ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //      avalon_anti_slave_0.read
		.av_readdata              (ifsr_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_address               (),                                                                                 //              (terminated)
		.av_write                 (),                                                                                 //              (terminated)
		.av_writedata             (),                                                                                 //              (terminated)
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_byteenable            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                      (clk_clk),                                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                                      //              (terminated)
		.av_read                  (),                                                                                      //              (terminated)
		.av_writedata             (),                                                                                      //              (terminated)
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_byteenable            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_ii_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                                //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.av_address              (nios_ii_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_ii_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_ii_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_ii_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_ii_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_ii_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_ii_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_ii_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_ii_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_ii_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_ii_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                                 //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                  //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                               //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                           //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                                 //          .ready
		.av_response             (),                                                                                       // (terminated)
		.av_writeresponserequest (1'b0),                                                                                   // (terminated)
		.av_writeresponsevalid   ()                                                                                        // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (71),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.PKT_BURST_TYPE_H          (68),
		.PKT_BURST_TYPE_L          (67),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_TRANS_EXCLUSIVE       (57),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (70),
		.PKT_DATA_SIDEBAND_L       (70),
		.PKT_QOS_H                 (72),
		.PKT_QOS_L                 (72),
		.PKT_ADDR_SIDEBAND_H       (69),
		.PKT_ADDR_SIDEBAND_L       (69),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_ii_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                         //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.av_address              (nios_ii_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios_ii_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios_ii_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios_ii_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios_ii_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios_ii_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios_ii_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios_ii_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios_ii_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios_ii_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios_ii_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                       //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                      //          .ready
		.av_response             (),                                                                                // (terminated)
		.av_writeresponserequest (1'b0),                                                                            // (terminated)
		.av_writeresponsevalid   ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                       //                .channel
		.rf_sink_ready           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                //                .channel
		.rf_sink_ready           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                       //     (terminated)
		.m0_writeresponserequest (),                                                                            //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                         //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                               //                .channel
		.rf_sink_ready           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                                    //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                                 //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (71),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (51),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (52),
		.PKT_TRANS_POSTED          (53),
		.PKT_TRANS_WRITE           (54),
		.PKT_TRANS_READ            (55),
		.PKT_TRANS_LOCK            (56),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (73),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (63),
		.PKT_BURSTWRAP_L           (61),
		.PKT_BYTE_CNT_H            (60),
		.PKT_BYTE_CNT_L            (58),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (66),
		.PKT_BURST_SIZE_L          (64),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                 //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	SOC_addr_router addr_router (
		.sink_ready         (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_ii_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_src_valid),                                                                  //          .valid
		.src_data           (addr_router_src_data),                                                                   //          .data
		.src_channel        (addr_router_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                             //          .endofpacket
	);

	SOC_addr_router_001 addr_router_001 (
		.sink_ready         (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_ii_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                       //          .valid
		.src_data           (addr_router_001_src_data),                                                        //          .data
		.src_channel        (addr_router_001_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                  //          .endofpacket
	);

	SOC_id_router id_router (
		.sink_ready         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios_ii_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_src_valid),                                                                  //          .valid
		.src_data           (id_router_src_data),                                                                   //          .data
		.src_channel        (id_router_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                             //          .endofpacket
	);

	SOC_id_router id_router_001 (
		.sink_ready         (ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                           //       src.ready
		.src_valid          (id_router_001_src_valid),                                           //          .valid
		.src_data           (id_router_001_src_data),                                            //          .data
		.src_channel        (id_router_001_src_channel),                                         //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                   //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                      //          .endofpacket
	);

	SOC_id_router id_router_002 (
		.sink_ready         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ifsr_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                          //       src.ready
		.src_valid          (id_router_002_src_valid),                                                          //          .valid
		.src_data           (id_router_002_src_data),                                                           //          .data
		.src_channel        (id_router_002_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                     //          .endofpacket
	);

	SOC_id_router_003 id_router_003 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                             //          .endofpacket
	);

	SOC_id_router_003 id_router_004 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                                               //          .valid
		.src_data           (id_router_004_src_data),                                                                //          .data
		.src_channel        (id_router_004_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                          //          .endofpacket
	);

	SOC_id_router_003 id_router_005 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                               //       src.ready
		.src_valid          (id_router_005_src_valid),                                               //          .valid
		.src_data           (id_router_005_src_data),                                                //          .data
		.src_channel        (id_router_005_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                          //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	SOC_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket)    //          .endofpacket
	);

	SOC_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //      src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	SOC_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	SOC_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SOC_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux_003 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	SOC_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	SOC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_ii_d_irq_irq)               //    sender.irq
	);

endmodule
